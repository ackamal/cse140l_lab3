// traffic light controller shell -- fill in the guts
// CSE140L  Summer II  2019
module traffic_light_controller(
  input clk,                          // 
        reset,						  // should force to all-red state
        ew_left_sensor,
        ew_str_sensor,	
        ns_sensor,
output logic[1:0] ew_left_light,     
			      ew_str_light,	
			      ns_light);



endmodule 